LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.math_real.ceil;

PACKAGE general_package IS
    -- DATA FORMAT
    CONSTANT N_BITS : INTEGER := 16;
    CONSTANT N_FLOAT : INTEGER := 0;

    -- ARCHITECTURE PARAMETERS
    CONSTANT N_UNITS : INTEGER := 32; -- MUST BE A POWER OF TWO
    CONSTANT N_PARALL : INTEGER := 4; -- MUST BE A POWER OF TWO LESS THAN N_UNITS
    CONSTANT DEPTH : INTEGER := INTEGER(ceil(real(N_UNITS/N_PARALL)));

    -- BUSES
    TYPE K_BUS IS ARRAY (N_PARALL - 1 DOWNTO 0) OF STD_LOGIC_VECTOR (N_BITS - 1 DOWNTO 0);
    TYPE N_BUS IS ARRAY (N_UNITS - 1 DOWNTO 0) OF STD_LOGIC_VECTOR (N_BITS - 1 DOWNTO 0);
    TYPE NK_BUS IS ARRAY (DEPTH - 1 DOWNTO 0) OF K_BUS;
END PACKAGE;